`define ADDR_WIDTH 8
`define DATA_WIDTH 32
`define MEM_DEPTH 256
`define STRB_WIDTH 4