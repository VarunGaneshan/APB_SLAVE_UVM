class apb_passive_monitor extends uvm_monitor;
  `uvm_component_utils(apb_passive_monitor)
  
  virtual apb_if vif;
  uvm_analysis_port#(apb_sequence_item) mon_port;
  apb_sequence_item mon_trans;
    
  function new(string name="apb_passive_monitor", uvm_component parent=null);
    super.new(name, parent);
    mon_port = new("mon_port", this);
  endfunction
    
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if(!uvm_config_db#(virtual apb_if)::get(this, "", "vif", vif)) begin
      `uvm_fatal("NOVIF", "No virtual interface found");
    end
  endfunction
  
  virtual task run_phase(uvm_phase phase);
    super.run_phase(phase);
    
    // Wait for reset deassertion
    @(posedge vif.presetn);
    `uvm_info(get_type_name(), $sformatf("[%0t] Reset De-asserted", $time), UVM_LOW)
    
    forever begin
      // Wait for valid APB transfer at clock edge
      @(posedge vif.pclk);
      
      if (vif.psel && vif.penable) begin
        // Capture inputs during ACCESS phase
        mon_trans = apb_sequence_item::type_id::create("mon_trans");
        
        // Wait one more clock to get registered outputs from DUT
        @(posedge vif.pclk);
        capture_outputs();
        
        // Send complete transaction to scoreboard and subscriber
        mon_port.write(mon_trans);
        
        `uvm_info(get_type_name(), 
                  $sformatf("[%0t] Captured Transaction: ADDR=0x%0h, WRITE=%0b, WDATA=0x%0h, STRB=0x%0h, RDATA=0x%0h, READY=%0b, SLVERR=%0b", 
                           $time,
                           mon_trans.paddr,
                           mon_trans.pwrite,
                           mon_trans.pwdata,
                           mon_trans.pstrb,
                           mon_trans.prdata, 
                           mon_trans.pready,
                           mon_trans.pslverr), 
                  UVM_MEDIUM)
      end
    end
  endtask             
         
  // Capture output signals after registered outputs update
  virtual task capture_outputs();
    mon_trans.prdata  = vif.prdata;
    mon_trans.pready  = vif.pready;
    mon_trans.pslverr = vif.pslverr;
  endtask
  
endclass
